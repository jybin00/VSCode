`include "TPMEM_16x16.v"

module 2D_DCT();


endmodule