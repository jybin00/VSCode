`include "rythm.v"
`timescale 1us/1us

module rtb;

menu1,