module tpmem_st2_opt
#( parameter BW = 12 )
// 입력 데이터, enable 신호, 입력 클럭, 입력 리셋, 출력 데이ㅓㅌ, 출력 enable 신호
(  input        [16*BW-1:0]	i_data,
   input	   	            i_enable,
   input 	   	            i_clk,
   input	   	            i_Reset,
   output reg   [16*BW-1:0] o_data,
   output reg	            o_en
);

// counter <= 입출력할 때 사용하려고 선언함.
reg [5-1:0]         counter;
reg [154-1:0] a0;
reg [148-1:0] a1;
reg [142-1:0] a2;
reg [140-1:0] a3;
reg [137-1:0] a4;
reg [133-1:0] a5;
reg [129-1:0] a6;
reg [130-1:0] a7;
reg [125-1:0] a8;
reg [123-1:0] a9;
reg [121-1:0] a10;
reg [122-1:0] a11;
reg [119-1:0] a12;
reg [120-1:0] a13;
reg [116-1:0] a14;
reg [116-1:0] a15;
// Data 출력을 위한 reg
reg [16*BW-1:0]     data_out;

// col은 말 그대로 column. 
wire [16*BW-1:0]    col     [16-1:0];
wire [4-1:0]        index = counter[4-1:0] ;

// Data 츌력 위한 wire
wire [16*BW-1:0]    w_data;
wire	            w_en;

wire signed [12-1:0] Xk_0 = i_data[15*12 +: 12];
wire signed [12-1:0] Xk_1 = i_data[14*12 +: 12];
wire signed [12-1:0] Xk_2 = i_data[13*12 +: 12];
wire signed [12-1:0] Xk_3 = i_data[12*12 +: 12];
wire signed [12-1:0] Xk_4 = i_data[11*12 +: 12];
wire signed [12-1:0] Xk_5 = i_data[10*12 +: 12];
wire signed [12-1:0] Xk_6 = i_data[ 9*12 +: 12];
wire signed [12-1:0] Xk_7 = i_data[ 8*12 +: 12];
wire signed [12-1:0] Xk_8 = i_data[ 7*12 +: 12];
wire signed [12-1:0] Xk_9 = i_data[ 6*12 +: 12];
wire signed [12-1:0] Xk_10 = i_data[ 5*12 +: 12];
wire signed [12-1:0] Xk_11 = i_data[ 4*12 +: 12];
wire signed [12-1:0] Xk_12 = i_data[ 3*12 +: 12];
wire signed [12-1:0] Xk_13 = i_data[ 2*12 +: 12];
wire signed [12-1:0] Xk_14 = i_data[ 1*12 +: 12];
wire signed [12-1:0] Xk_15 = i_data[ 0*12 +: 12];


always@(posedge i_clk) begin
    if(~i_Reset) begin
        // counter, o_data, o_en 초기화
        counter <= 5'b0;
        o_data  <= {BW{16'b0}};
        o_en    <= 1'b0; 
    end
    else begin
        // o_data에는 w_data를, o_en에는 w_en을 대입
        o_data  <= w_data ;
        o_en    <= w_en ;
        if(i_enable) 
            // input이 enable일 때. counter를 1씩 증가시킴.
            counter     <= counter + 5'b1;
        else begin  
            // input이 enable이 아니면서, counter[4]가 1일 때.  
            // 카운터가 증가하면 index도 1씩 증가함.
            if(counter[4]==1'b1) counter <= counter + 5'b1;
    	    else counter <= counter ;
    	end
    end
end

always@(posedge i_clk) begin
    if(~i_Reset) begin
        // array 초기화
        a0  <= {154'b0};
        a1  <= {148'b0};
        a2  <= {142'b0};
        a3  <= {140'b0};
        a4  <= {137'b0};
        a5  <= {133'b0};
        a6  <= {129'b0};
        a7  <= {130'b0};
        a8  <= {125'b0};
        a9  <= {123'b0};
        a10 <= {121'b0};
        a11 <= {122'b0};
        a12 <= {119'b0};
        a13 <= {120'b0};
        a14 <= {116'b0};
        a15 <= {116'b0};
    end
    else begin
        if(i_enable) begin
            // reset 아니고 enable일 때, array에 i_data를 대입함.
            case(index)
                4'b0000: a0  <= {Xk_0,        Xk_1,         Xk_2,        Xk_3,         Xk_4[10-1:0], Xk_5[10-1:0],Xk_6[10-1:0],Xk_7[9-1:0], Xk_8[9-1:0], Xk_9[9-1:0], Xk_10[8-1:0], Xk_11[8-1:0], Xk_12[8-1:0], Xk_13[9-1:0], Xk_14[8-1:0], Xk_15[8-1:0]};
                4'b0001: a1  <= {Xk_0,        Xk_1,         Xk_2,        Xk_3[10-1:0], Xk_4[10-1:0], Xk_5[9-1:0], Xk_6[9-1:0], Xk_7[9-1:0], Xk_8[9-1:0], Xk_9[8-1:0], Xk_10[8-1:0], Xk_11[8-1:0], Xk_12[8-1:0], Xk_13[8-1:0], Xk_14[8-1:0], Xk_15[8-1:0]};
                4'b0010: a2  <= {Xk_0,        Xk_1[10-1:0], Xk_2[10-1:0],Xk_3[10-1:0], Xk_4[10-1:0], Xk_5[9-1:0], Xk_6[9-1:0], Xk_7[8-1:0], Xk_8[8-1:0], Xk_9[8-1:0], Xk_10[8-1:0], Xk_11[8-1:0], Xk_12[8-1:0], Xk_13[8-1:0], Xk_14[8-1:0], Xk_15[8-1:0]};
                4'b0011: a3  <= {Xk_0[10-1:0],Xk_1[10-1:0], Xk_2[10-1:0],Xk_3[10-1:0], Xk_4[10-1:0], Xk_5[9-1:0], Xk_6[9-1:0], Xk_7[8-1:0], Xk_8[8-1:0], Xk_9[8-1:0], Xk_10[8-1:0], Xk_11[8-1:0], Xk_12[8-1:0], Xk_13[8-1:0], Xk_14[8-1:0], Xk_15[8-1:0]};
                4'b0100: a4  <= {Xk_0[10-1:0],Xk_1[10-1:0], Xk_2[10-1:0],Xk_3[9-1:0],  Xk_4[9-1:0],  Xk_5[9-1:0], Xk_6[8-1:0], Xk_7[8-1:0], Xk_8[8-1:0], Xk_9[8-1:0], Xk_10[8-1:0], Xk_11[8-1:0], Xk_12[8-1:0], Xk_13[8-1:0], Xk_14[8-1:0], Xk_15[8-1:0]};
                4'b0101: a5  <= {Xk_0[10-1:0],Xk_1[10-1:0], Xk_2[9-1:0], Xk_3[9-1:0],  Xk_4[9-1:0],  Xk_5[9-1:0], Xk_6[8-1:0], Xk_7[8-1:0], Xk_8[8-1:0], Xk_9[8-1:0], Xk_10[8-1:0], Xk_11[8-1:0], Xk_12[8-1:0], Xk_13[8-1:0], Xk_14[8-1:0], Xk_15[8-1:0]};
                4'b0110: a6  <= {Xk_0[10-1:0],Xk_1[10-1:0], Xk_2[9-1:0], Xk_3[9-1:0],  Xk_4[9-1:0],  Xk_5[8-1:0], Xk_6[8-1:0], Xk_7[8-1:0], Xk_8[8-1:0], Xk_9[8-1:0], Xk_10[7-1:0], Xk_11[7-1:0], Xk_12[7-1:0], Xk_13[7-1:0], Xk_14[7-1:0], Xk_15[7-1:0]};
                4'b0111: a7  <= {Xk_0        ,Xk_1[10-1:0], Xk_2[9-1:0], Xk_3[9-1:0],  Xk_4[8-1:0],  Xk_5[8-1:0], Xk_6[8-1:0], Xk_7[8-1:0], Xk_8[8-1:0], Xk_9[8-1:0], Xk_10[7-1:0], Xk_11[7-1:0], Xk_12[7-1:0], Xk_13[7-1:0], Xk_14[7-1:0], Xk_15[7-1:0]};
                4'b1000: a8  <= {Xk_0[10-1:0],Xk_1[9 -1:0], Xk_2[8-1:0], Xk_3[8-1:0],  Xk_4[8-1:0],  Xk_5[8-1:0], Xk_6[8-1:0], Xk_7[8-1:0], Xk_8[8-1:0], Xk_9[8-1:0], Xk_10[7-1:0], Xk_11[7-1:0], Xk_12[7-1:0], Xk_13[7-1:0], Xk_14[7-1:0], Xk_15[7-1:0]};
                4'b1001: a9  <= {Xk_0[9 -1:0], Xk_1[8-1:0], Xk_2[8-1:0], Xk_3[8-1:0],  Xk_4[8-1:0],  Xk_5[8-1:0], Xk_6[8-1:0], Xk_7[8-1:0], Xk_8[8-1:0], Xk_9[8-1:0], Xk_10[7-1:0], Xk_11[7-1:0], Xk_12[7-1:0], Xk_13[7-1:0], Xk_14[7-1:0], Xk_15[7-1:0]};
                4'b1010: a10 <= {Xk_0[9 -1:0], Xk_1[8-1:0], Xk_2[8-1:0], Xk_3[9-1:0],  Xk_4[8-1:0],  Xk_5[8-1:0], Xk_6[8-1:0], Xk_7[7-1:0], Xk_8[7-1:0], Xk_9[7-1:0], Xk_10[7-1:0], Xk_11[7-1:0], Xk_12[7-1:0], Xk_13[7-1:0], Xk_14[7-1:0], Xk_15[7-1:0]};
                4'b1011: a11 <= {Xk_0[9 -1:0], Xk_1[8-1:0], Xk_2[9-1:0], Xk_3[8-1:0],  Xk_4[9-1:0],  Xk_5[8-1:0], Xk_6[8-1:0], Xk_7[7-1:0], Xk_8[7-1:0], Xk_9[7-1:0], Xk_10[7-1:0], Xk_11[7-1:0], Xk_12[7-1:0], Xk_13[7-1:0], Xk_14[7-1:0], Xk_15[7-1:0]};
                4'b1100: a12 <= {Xk_0[8 -1:0], Xk_1[8-1:0], Xk_2[8-1:0], Xk_3[8-1:0],  Xk_4[8-1:0],  Xk_5[8-1:0], Xk_6[8-1:0], Xk_7[7-1:0], Xk_8[7-1:0], Xk_9[7-1:0], Xk_10[7-1:0], Xk_11[7-1:0], Xk_12[7-1:0], Xk_13[7-1:0], Xk_14[7-1:0], Xk_15[7-1:0]};
                4'b1101: a13 <= {Xk_0[8 -1:0], Xk_1[8-1:0], Xk_2[8-1:0], Xk_3[8-1:0],  Xk_4[8-1:0],  Xk_5[8-1:0], Xk_6[8-1:0], Xk_7[7-1:0], Xk_8[7-1:0], Xk_9[8-1:0], Xk_10[7-1:0], Xk_11[7-1:0], Xk_12[7-1:0], Xk_13[7-1:0], Xk_14[7-1:0], Xk_15[7-1:0]};
                4'b1110: a14 <= {Xk_0[8 -1:0], Xk_1[8-1:0], Xk_2[8-1:0], Xk_3[8-1:0],  Xk_4[7-1:0],  Xk_5[7-1:0], Xk_6[7-1:0], Xk_7[7-1:0], Xk_8[7-1:0], Xk_9[7-1:0], Xk_10[7-1:0], Xk_11[7-1:0], Xk_12[7-1:0], Xk_13[7-1:0], Xk_14[7-1:0], Xk_15[7-1:0]};
                4'b1111: a15 <= {Xk_0[8 -1:0], Xk_1[8-1:0], Xk_2[8-1:0], Xk_3[8-1:0],  Xk_4[7-1:0],  Xk_5[7-1:0], Xk_6[7-1:0], Xk_7[7-1:0], Xk_8[7-1:0], Xk_9[7-1:0], Xk_10[7-1:0], Xk_11[7-1:0], Xk_12[7-1:0], Xk_13[7-1:0], Xk_14[7-1:0], Xk_15[7-1:0]};
            endcase
            //array[index] <= i_data ;
        end
    end
end

assign col[ 0] = {{a0[154-1:142]},             {a1[16*BW-1:15*BW]},{a2[16*BW-1:15*BW]},{a3[16*BW-1:15*BW]},{a4[16*BW-1:15*BW]},{a5[16*BW-1:15*BW]},{a6[16*BW-1:15*BW]},{a7[16*BW-1:15*BW]},{a8[16*BW-1:15*BW]},{a9[16*BW-1:15*BW]},{a10[16*BW-1:15*BW]},{a11[16*BW-1:15*BW]},{a12[16*BW-1:15*BW]},{a13[16*BW-1:15*BW]},{a14[16*BW-1:15*BW]},{a15[16*BW-1:15*BW]}} ; 
assign col[ 1] = {{a0[142-1:130]},             {a1[15*BW-1:14*BW]},{a2[15*BW-1:14*BW]},{a3[15*BW-1:14*BW]},{a4[15*BW-1:14*BW]},{a5[15*BW-1:14*BW]},{a6[15*BW-1:14*BW]},{a7[15*BW-1:14*BW]},{a8[15*BW-1:14*BW]},{a9[15*BW-1:14*BW]},{a10[15*BW-1:14*BW]},{a11[15*BW-1:14*BW]},{a12[15*BW-1:14*BW]},{a13[15*BW-1:14*BW]},{a14[15*BW-1:14*BW]},{a15[15*BW-1:14*BW]}} ; 
assign col[ 2] = {{a0[130-1:118]},             {a1[14*BW-1:13*BW]},{a2[14*BW-1:13*BW]},{a3[14*BW-1:13*BW]},{a4[14*BW-1:13*BW]},{a5[14*BW-1:13*BW]},{a6[14*BW-1:13*BW]},{a7[14*BW-1:13*BW]},{a8[14*BW-1:13*BW]},{a9[14*BW-1:13*BW]},{a10[14*BW-1:13*BW]},{a11[14*BW-1:13*BW]},{a12[14*BW-1:13*BW]},{a13[14*BW-1:13*BW]},{a14[14*BW-1:13*BW]},{a15[14*BW-1:13*BW]}} ; 
assign col[ 3] = {{a0[118-1:106]},             {a1[13*BW-1:12*BW]},{a2[13*BW-1:12*BW]},{a3[13*BW-1:12*BW]},{a4[13*BW-1:12*BW]},{a5[13*BW-1:12*BW]},{a6[13*BW-1:12*BW]},{a7[13*BW-1:12*BW]},{a8[13*BW-1:12*BW]},{a9[13*BW-1:12*BW]},{a10[13*BW-1:12*BW]},{a11[13*BW-1:12*BW]},{a12[13*BW-1:12*BW]},{a13[13*BW-1:12*BW]},{a14[13*BW-1:12*BW]},{a15[13*BW-1:12*BW]}} ; 
assign col[ 4] = {{{2{a0[105]}},a0[106-1: 96]},{a1[12*BW-1:11*BW]},{a2[12*BW-1:11*BW]},{a3[12*BW-1:11*BW]},{a4[12*BW-1:11*BW]},{a5[12*BW-1:11*BW]},{a6[12*BW-1:11*BW]},{a7[12*BW-1:11*BW]},{a8[12*BW-1:11*BW]},{a9[12*BW-1:11*BW]},{a10[12*BW-1:11*BW]},{a11[12*BW-1:11*BW]},{a12[12*BW-1:11*BW]},{a13[12*BW-1:11*BW]},{a14[12*BW-1:11*BW]},{a15[12*BW-1:11*BW]}} ; 
assign col[ 5] = {{a0[ 96-1: 86]},             {a1[11*BW-1:10*BW]},{a2[11*BW-1:10*BW]},{a3[11*BW-1:10*BW]},{a4[11*BW-1:10*BW]},{a5[11*BW-1:10*BW]},{a6[11*BW-1:10*BW]},{a7[11*BW-1:10*BW]},{a8[11*BW-1:10*BW]},{a9[11*BW-1:10*BW]},{a10[11*BW-1:10*BW]},{a11[11*BW-1:10*BW]},{a12[11*BW-1:10*BW]},{a13[11*BW-1:10*BW]},{a14[11*BW-1:10*BW]},{a15[11*BW-1:10*BW]}} ; 
assign col[ 6] = {{a0[ 86-1: 76]},             {a1[10*BW-1: 9*BW]},{a2[10*BW-1: 9*BW]},{a3[10*BW-1: 9*BW]},{a4[10*BW-1: 9*BW]},{a5[10*BW-1: 9*BW]},{a6[10*BW-1: 9*BW]},{a7[10*BW-1: 9*BW]},{a8[10*BW-1: 9*BW]},{a9[10*BW-1: 9*BW]},{a10[10*BW-1: 9*BW]},{a11[10*BW-1: 9*BW]},{a12[10*BW-1: 9*BW]},{a13[10*BW-1: 9*BW]},{a14[10*BW-1: 9*BW]},{a15[10*BW-1: 9*BW]}} ;
assign col[ 7] = {{a0[ 76-1: 67]},             {a1[ 9*BW-1: 8*BW]},{a2[ 9*BW-1: 8*BW]},{a3[ 9*BW-1: 8*BW]},{a4[ 9*BW-1: 8*BW]},{a5[ 9*BW-1: 8*BW]},{a6[ 9*BW-1: 8*BW]},{a7[ 9*BW-1: 8*BW]},{a8[ 9*BW-1: 8*BW]},{a9[ 9*BW-1: 8*BW]},{a10[ 9*BW-1: 8*BW]},{a11[ 9*BW-1: 8*BW]},{a12[ 9*BW-1: 8*BW]},{a13[ 9*BW-1: 8*BW]},{a14[ 9*BW-1: 8*BW]},{a15[ 9*BW-1: 8*BW]}} ;

assign col[ 8] = {{a0[067-1:058]},             {a1[ 8*BW-1: 7*BW]},{a2[ 8*BW-1: 7*BW]},{a3[ 8*BW-1: 7*BW]},{a4[ 8*BW-1: 7*BW]},{a5[ 8*BW-1: 7*BW]},{a6[ 8*BW-1: 7*BW]},{a7[ 8*BW-1: 7*BW]},{a8[ 8*BW-1: 7*BW]},{a9[ 8*BW-1: 7*BW]},{a10[ 8*BW-1: 7*BW]},{a11[ 8*BW-1: 7*BW]},{a12[ 8*BW-1: 7*BW]},{a13[ 8*BW-1: 7*BW]},{a14[ 8*BW-1: 7*BW]},{a15[ 8*BW-1: 7*BW]}} ; 
assign col[ 9] = {{a0[058-1:049]},             {a1[ 7*BW-1: 6*BW]},{a2[ 7*BW-1: 6*BW]},{a3[ 7*BW-1: 6*BW]},{a4[ 7*BW-1: 6*BW]},{a5[ 7*BW-1: 6*BW]},{a6[ 7*BW-1: 6*BW]},{a7[ 7*BW-1: 6*BW]},{a8[ 7*BW-1: 6*BW]},{a9[ 7*BW-1: 6*BW]},{a10[ 7*BW-1: 6*BW]},{a11[ 7*BW-1: 6*BW]},{a12[ 7*BW-1: 6*BW]},{a13[ 7*BW-1: 6*BW]},{a14[ 7*BW-1: 6*BW]},{a15[ 7*BW-1: 6*BW]}} ; 
assign col[10] = {{a0[049-1:041]},             {a1[ 6*BW-1: 5*BW]},{a2[ 6*BW-1: 5*BW]},{a3[ 6*BW-1: 5*BW]},{a4[ 6*BW-1: 5*BW]},{a5[ 6*BW-1: 5*BW]},{a6[ 6*BW-1: 5*BW]},{a7[ 6*BW-1: 5*BW]},{a8[ 6*BW-1: 5*BW]},{a9[ 6*BW-1: 5*BW]},{a10[ 6*BW-1: 5*BW]},{a11[ 6*BW-1: 5*BW]},{a12[ 6*BW-1: 5*BW]},{a13[ 6*BW-1: 5*BW]},{a14[ 6*BW-1: 5*BW]},{a15[ 6*BW-1: 5*BW]}} ; 
assign col[11] = {{a0[041-1:033]},             {a1[ 5*BW-1: 4*BW]},{a2[ 5*BW-1: 4*BW]},{a3[ 5*BW-1: 4*BW]},{a4[ 5*BW-1: 4*BW]},{a5[ 5*BW-1: 4*BW]},{a6[ 5*BW-1: 4*BW]},{a7[ 5*BW-1: 4*BW]},{a8[ 5*BW-1: 4*BW]},{a9[ 5*BW-1: 4*BW]},{a10[ 5*BW-1: 4*BW]},{a11[ 5*BW-1: 4*BW]},{a12[ 5*BW-1: 4*BW]},{a13[ 5*BW-1: 4*BW]},{a14[ 5*BW-1: 4*BW]},{a15[ 5*BW-1: 4*BW]}} ; 
assign col[12] = {{a0[033-1:025]},             {a1[ 4*BW-1: 3*BW]},{a2[ 4*BW-1: 3*BW]},{a3[ 4*BW-1: 3*BW]},{a4[ 4*BW-1: 3*BW]},{a5[ 4*BW-1: 3*BW]},{a6[ 4*BW-1: 3*BW]},{a7[ 4*BW-1: 3*BW]},{a8[ 4*BW-1: 3*BW]},{a9[ 4*BW-1: 3*BW]},{a10[ 4*BW-1: 3*BW]},{a11[ 4*BW-1: 3*BW]},{a12[ 4*BW-1: 3*BW]},{a13[ 4*BW-1: 3*BW]},{a14[ 4*BW-1: 3*BW]},{a15[ 4*BW-1: 3*BW]}} ; 
assign col[13] = {{a0[025-1:016]},             {a1[ 3*BW-1: 2*BW]},{a2[ 3*BW-1: 2*BW]},{a3[ 3*BW-1: 2*BW]},{a4[ 3*BW-1: 2*BW]},{a5[ 3*BW-1: 2*BW]},{a6[ 3*BW-1: 2*BW]},{a7[ 3*BW-1: 2*BW]},{a8[ 3*BW-1: 2*BW]},{a9[ 3*BW-1: 2*BW]},{a10[ 3*BW-1: 2*BW]},{a11[ 3*BW-1: 2*BW]},{a12[ 3*BW-1: 2*BW]},{a13[ 3*BW-1: 2*BW]},{a14[ 3*BW-1: 2*BW]},{a15[ 3*BW-1: 2*BW]}} ; 
assign col[14] = {{a0[016-1:008]},             {a1[ 2*BW-1: 1*BW]},{a2[ 2*BW-1: 1*BW]},{a3[ 2*BW-1: 1*BW]},{a4[ 2*BW-1: 1*BW]},{a5[ 2*BW-1: 1*BW]},{a6[ 2*BW-1: 1*BW]},{a7[ 2*BW-1: 1*BW]},{a8[ 2*BW-1: 1*BW]},{a9[ 2*BW-1: 1*BW]},{a10[ 2*BW-1: 1*BW]},{a11[ 2*BW-1: 1*BW]},{a12[ 2*BW-1: 1*BW]},{a13[ 2*BW-1: 1*BW]},{a14[ 2*BW-1: 1*BW]},{a15[ 2*BW-1: 1*BW]}} ;
assign col[15] = {{a0[008-1:000]},             {a1[ 1*BW-1: 0*BW]},{a2[ 1*BW-1: 0*BW]},{a3[ 1*BW-1: 0*BW]},{a4[ 1*BW-1: 0*BW]},{a5[ 1*BW-1: 0*BW]},{a6[ 1*BW-1: 0*BW]},{a7[ 1*BW-1: 0*BW]},{a8[ 1*BW-1: 0*BW]},{a9[ 1*BW-1: 0*BW]},{a10[ 1*BW-1: 0*BW]},{a11[ 1*BW-1: 0*BW]},{a12[ 1*BW-1: 0*BW]},{a13[ 1*BW-1: 0*BW]},{a14[ 1*BW-1: 0*BW]},{a15[ 1*BW-1: 0*BW]}} ;
always@(*) begin
    if(counter[4]==1'b1) data_out = col[index] ;
    else data_out = {BW{16'b0}}; 
end

assign w_en = counter[4] ;
assign w_data = data_out ; 

endmodule
