
module direct_filt(direct_out, direct_in, clk, rstn, c0, c1, c2, c3, c4);
    output signed[22-1:0] direct_out;
    input signed [12-1:0] direct_in;
    input clk, rstn;
    input signed[12-1:0] c0, c1, c2, c3, c4;



endmodule